`timescale 1ns / 1ps

module SDLC_result(
    input  [14:0] R1, R2, R3, R4,
    output [15:0] S
);

    // Verilog�� + �����ڴ� �ջ� ����� ����� ��Ʈ ������ �ڵ� Ȯ���մϴ�.
    // 15��Ʈ ���� 4���� ���ϸ� ����� �ִ� 17��Ʈ�� �� �� �����Ƿ�,
    // �׿� ���� �߰� ����� ���� ����� �����ϴ� ���� �����ϴ�.
    wire [16:0] temp_sum;
    
    // �� ���� �Է��� �� ���� ���մϴ�.
    // �ռ� ������ �� �ڵ带 ���� ���������� ȿ������ ���� Ʈ�� ������ �����մϴ�.
    assign temp_sum = R1 + R2 + R3 + R4;

    // ���� ��� S�� 16��Ʈ�̹Ƿ�, ��� ����� ���� 16��Ʈ�� �Ҵ��մϴ�.
    // ���� 17��Ʈ ��ü ����� �ʿ��ϴٸ� output S�� [16:0]���� �����ؾ� �մϴ�.
    assign S = temp_sum[15:0];

endmodule